

black   := "000";
blue    := "001";
green   := "010";
cyan    := "011";
red     := "100";
magenta := "101";
yellow  := "110";
white   := "111";
